
library ieee;
use ieee.std_logic_1164.all;

library work;
use work.lab4_pck.all;

library work;
use work.all;
use work.lab4_tb_pck.all;

entity tb_lab4 is
  
  -- empty signal list
end tb_lab4;
